library verilog;
use verilog.vl_types.all;
entity mean_filter_tb is
end mean_filter_tb;
